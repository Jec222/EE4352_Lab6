module and1 (z,a,b);
output z;
input a,b;
assign  z= a & b;
endmodule